library verilog;
use verilog.vl_types.all;
entity StoreSize_vlg_vec_tst is
end StoreSize_vlg_vec_tst;
