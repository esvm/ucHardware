library verilog;
use verilog.vl_types.all;
entity Div_vlg_vec_tst is
end Div_vlg_vec_tst;
