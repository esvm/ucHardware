library verilog;
use verilog.vl_types.all;
entity LoadSize is
    port(
        LSControl       : in     vl_logic_vector(1 downto 0);
        Data            : in     vl_logic_vector(31 downto 0);
        \out\           : out    vl_logic_vector(31 downto 0)
    );
end LoadSize;
