library verilog;
use verilog.vl_types.all;
entity ShiftLeft16_vlg_vec_tst is
end ShiftLeft16_vlg_vec_tst;
