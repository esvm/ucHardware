library verilog;
use verilog.vl_types.all;
entity LoadSize_vlg_vec_tst is
end LoadSize_vlg_vec_tst;
